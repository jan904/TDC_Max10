-- State machine for handling the signal detection. Once a input signal is detected,
-- signal_running is set to '1' to lock the FFs of the delay line. Then wrt is set to '1'
-- to write the signal to the FIFO. Once the signal is written, reset is set to '1' to reset the delay line. 

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY detect_signal IS
    GENERIC (
        stages : INTEGER := 124;                    -- Number of bins in the delay line
        n_output_bits : INTEGER := 8                -- Number of bits for fine timestamp
    );
    PORT (
        clock : IN STD_LOGIC;                       -- Clock 
        start : IN STD_LOGIC;                       -- Reset signal after start of the FPGA. Generated by handle_start
        signal_in : IN STD_LOGIC;                   -- Input signal which is to be detected
        written : IN STD_LOGIC;                     -- Signal to indicate that the output of this channel has been written to the FIFO
        signal_running : OUT STD_LOGIC;             -- Signal to indicate that the delay chain is busy with a signal
        reset : OUT STD_LOGIC;                      -- Reset signal after signal has been processed
        wrt : OUT STD_LOGIC                         -- Write enable: Indicates that the output of this channel is ready to be written to the FIFO
    );
END ENTITY detect_signal;


ARCHITECTURE fsm OF detect_signal IS

    -- Define the states of the FSM
    TYPE stype IS (IDLE, DETECT_START, WRITE_FIFO, RST);
    SIGNAL state, next_state : stype;

    -- Signals used to store the values of the signals
    SIGNAL reset_reg, reset_next : STD_LOGIC;
    SIGNAL signal_running_reg, signal_running_next : STD_LOGIC;
    SIGNAL wrt_reg, wrt_next : STD_LOGIC;
    SIGNAL count, count_reg, count_next : INTEGER range 0 to 4;

BEGIN
    -- FSM core
    PROCESS(clock)
    BEGIN
        IF rising_edge(clock) THEN
            -- Reset at start 
            IF start = '1' THEN
                state <= IDLE;
                signal_running_reg <= '0';
                reset_reg <= '0';
                wrt_reg <= '0';
                count <= 0;

            -- Update signals
            ELSE
                signal_running_reg <= signal_running_next;
                reset_reg <= reset_next;
                wrt_reg <= wrt_next;
                state <= next_state;
                count <= count_next;
            END IF;
        END IF;
    END PROCESS;

    -- FSM logic
    PROCESS (state, signal_running_reg, wrt_reg, reset_reg, signal_in, count, written)  
    BEGIN

        -- Default values
        next_state <= state;
        wrt_next <= wrt_reg;
        reset_next <= reset_reg;
        signal_running_next <= signal_running_reg;
        count_next <= count;

        CASE state IS
            WHEN IDLE =>
                -- Start signal detection
                IF signal_in = '1' THEN
                    next_state <= DETECT_START;
                ELSE
                    next_state <= IDLE;
                END IF;
                
            WHEN DETECT_START =>
                -- Update signal_running to lock the delay line
                signal_running_next <= '1';
                next_state <= WRITE_FIFO;

            WHEN WRITE_FIFO =>
                -- Wait for three cycle for timing reasons. For some reason, using 3 separate IFs is much more stable than using "count < 3" statement
                IF count = 0 THEN
                    count_next <= count + 1;
                    next_state <= WRITE_FIFO;

                ELSIF count = 1 THEN
                    count_next <= count + 1;
                    next_state <= WRITE_FIFO;

                ELSIF count = 2 THEN
                    count_next <= count + 1;
                    next_state <= WRITE_FIFO;

                -- Enable wrt
                ELSIF count = 3 THEN
                    wrt_next <= '1';
                    count_next <= count + 1;
                    next_state <= WRITE_FIFO;

                -- If signal has been written, go to reset
                ELSIF count = 4 THEN
                    IF written = '1' THEN
                        next_state <= RST;
                    ELSE
                        next_state <= WRITE_FIFO;
                    END IF;

                -- If illegal state for some reason, go to reset
                ELSE
                    next_state <= RST;
                END IF;

            WHEN RST =>
                -- Wait until input is '0'. Then set reset to '1' for one cycle and return to idle
                -- Reset_reg ensures that the reset signal is only set for one cycle and the process does not
                -- get stuck if signal_in switches to '1' again (If this happens, the delay line records max value which should actually not happen)
                IF signal_in = '0' or reset_reg = '1' THEN
                    IF reset_reg = '1' THEN
                        next_state <= IDLE;
                        signal_running_next <= '0';
                        reset_next <= '0';
                        count_next <= 0;
                    ELSIF reset_reg = '0' THEN
                        next_state <= RST;
                        reset_next <= '1';
                    END IF;
                ELSE 
                    next_state <= RST;
                END IF;

                -- Default values
                wrt_next <= '0';

            -- Catch illegal states
            WHEN OTHERS =>
                next_state <= IDLE;
        END CASE;
    END PROCESS;

    -- Output signals
    signal_running <= signal_running_reg;
    reset <= reset_reg;
    wrt <= wrt_reg;

END ARCHITECTURE fsm;


