-- ethernet_setup.vhd

-- Generated using ACDS version 23.1 993

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity ethernet_setup is
	port (
		altpll_0_areset_conduit_export              : in  std_logic                     := '0';             --         altpll_0_areset_conduit.export
		altpll_0_c2_clk                             : out std_logic;                                        --                     altpll_0_c2.clk
		altpll_0_locked_conduit_export              : out std_logic;                                        --         altpll_0_locked_conduit.export
		clk_clk                                     : in  std_logic                     := '0';             --                             clk.clk
		eth_tse_0_mac_misc_connection_ff_tx_crc_fwd : in  std_logic                     := '0';             --   eth_tse_0_mac_misc_connection.ff_tx_crc_fwd
		eth_tse_0_mac_misc_connection_ff_tx_septy   : out std_logic;                                        --                                .ff_tx_septy
		eth_tse_0_mac_misc_connection_tx_ff_uflow   : out std_logic;                                        --                                .tx_ff_uflow
		eth_tse_0_mac_misc_connection_ff_tx_a_full  : out std_logic;                                        --                                .ff_tx_a_full
		eth_tse_0_mac_misc_connection_ff_tx_a_empty : out std_logic;                                        --                                .ff_tx_a_empty
		eth_tse_0_mac_misc_connection_rx_err_stat   : out std_logic_vector(17 downto 0);                    --                                .rx_err_stat
		eth_tse_0_mac_misc_connection_rx_frm_type   : out std_logic_vector(3 downto 0);                     --                                .rx_frm_type
		eth_tse_0_mac_misc_connection_ff_rx_dsav    : out std_logic;                                        --                                .ff_rx_dsav
		eth_tse_0_mac_misc_connection_ff_rx_a_full  : out std_logic;                                        --                                .ff_rx_a_full
		eth_tse_0_mac_misc_connection_ff_rx_a_empty : out std_logic;                                        --                                .ff_rx_a_empty
		eth_tse_0_mac_rgmii_connection_rgmii_in     : in  std_logic_vector(3 downto 0)  := (others => '0'); --  eth_tse_0_mac_rgmii_connection.rgmii_in
		eth_tse_0_mac_rgmii_connection_rgmii_out    : out std_logic_vector(3 downto 0);                     --                                .rgmii_out
		eth_tse_0_mac_rgmii_connection_rx_control   : in  std_logic                     := '0';             --                                .rx_control
		eth_tse_0_mac_rgmii_connection_tx_control   : out std_logic;                                        --                                .tx_control
		eth_tse_0_mac_status_connection_set_10      : in  std_logic                     := '0';             -- eth_tse_0_mac_status_connection.set_10
		eth_tse_0_mac_status_connection_set_1000    : in  std_logic                     := '0';             --                                .set_1000
		eth_tse_0_mac_status_connection_eth_mode    : out std_logic;                                        --                                .eth_mode
		eth_tse_0_mac_status_connection_ena_10      : out std_logic;                                        --                                .ena_10
		eth_tse_0_receive_data                      : out std_logic_vector(31 downto 0);                    --               eth_tse_0_receive.data
		eth_tse_0_receive_endofpacket               : out std_logic;                                        --                                .endofpacket
		eth_tse_0_receive_error                     : out std_logic_vector(5 downto 0);                     --                                .error
		eth_tse_0_receive_empty                     : out std_logic_vector(1 downto 0);                     --                                .empty
		eth_tse_0_receive_ready                     : in  std_logic                     := '0';             --                                .ready
		eth_tse_0_receive_startofpacket             : out std_logic;                                        --                                .startofpacket
		eth_tse_0_receive_valid                     : out std_logic;                                        --                                .valid
		eth_tse_0_transmit_data                     : in  std_logic_vector(31 downto 0) := (others => '0'); --              eth_tse_0_transmit.data
		eth_tse_0_transmit_endofpacket              : in  std_logic                     := '0';             --                                .endofpacket
		eth_tse_0_transmit_error                    : in  std_logic                     := '0';             --                                .error
		eth_tse_0_transmit_empty                    : in  std_logic_vector(1 downto 0)  := (others => '0'); --                                .empty
		eth_tse_0_transmit_ready                    : out std_logic;                                        --                                .ready
		eth_tse_0_transmit_startofpacket            : in  std_logic                     := '0';             --                                .startofpacket
		eth_tse_0_transmit_valid                    : in  std_logic                     := '0';             --                                .valid
		reset_reset_n                               : in  std_logic                     := '0'              --                           reset.reset_n
	);
end entity ethernet_setup;

architecture rtl of ethernet_setup is
	component ethernet_setup_altpll_0 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			read               : in  std_logic                     := 'X';             -- read
			write              : in  std_logic                     := 'X';             -- write
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0                 : out std_logic;                                        -- clk
			c1                 : out std_logic;                                        -- clk
			c2                 : out std_logic;                                        -- clk
			areset             : in  std_logic                     := 'X';             -- export
			locked             : out std_logic;                                        -- export
			scandone           : out std_logic;                                        -- export
			scandataout        : out std_logic;                                        -- export
			c3                 : out std_logic;                                        -- clk
			c4                 : out std_logic;                                        -- clk
			phasedone          : out std_logic;                                        -- export
			phasecounterselect : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- export
			phaseupdown        : in  std_logic                     := 'X';             -- export
			phasestep          : in  std_logic                     := 'X';             -- export
			scanclk            : in  std_logic                     := 'X';             -- export
			scanclkena         : in  std_logic                     := 'X';             -- export
			scandata           : in  std_logic                     := 'X';             -- export
			configupdate       : in  std_logic                     := 'X'              -- export
		);
	end component ethernet_setup_altpll_0;

	component ethernet_setup_eth_tse_0 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset         : in  std_logic                     := 'X';             -- reset
			reg_addr      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			reg_data_out  : out std_logic_vector(31 downto 0);                    -- readdata
			reg_rd        : in  std_logic                     := 'X';             -- read
			reg_data_in   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			reg_wr        : in  std_logic                     := 'X';             -- write
			reg_busy      : out std_logic;                                        -- waitrequest
			tx_clk        : in  std_logic                     := 'X';             -- clk
			rx_clk        : in  std_logic                     := 'X';             -- clk
			set_10        : in  std_logic                     := 'X';             -- set_10
			set_1000      : in  std_logic                     := 'X';             -- set_1000
			eth_mode      : out std_logic;                                        -- eth_mode
			ena_10        : out std_logic;                                        -- ena_10
			rgmii_in      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- rgmii_in
			rgmii_out     : out std_logic_vector(3 downto 0);                     -- rgmii_out
			rx_control    : in  std_logic                     := 'X';             -- rx_control
			tx_control    : out std_logic;                                        -- tx_control
			ff_rx_clk     : in  std_logic                     := 'X';             -- clk
			ff_tx_clk     : in  std_logic                     := 'X';             -- clk
			ff_rx_data    : out std_logic_vector(31 downto 0);                    -- data
			ff_rx_eop     : out std_logic;                                        -- endofpacket
			rx_err        : out std_logic_vector(5 downto 0);                     -- error
			ff_rx_mod     : out std_logic_vector(1 downto 0);                     -- empty
			ff_rx_rdy     : in  std_logic                     := 'X';             -- ready
			ff_rx_sop     : out std_logic;                                        -- startofpacket
			ff_rx_dval    : out std_logic;                                        -- valid
			ff_tx_data    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			ff_tx_eop     : in  std_logic                     := 'X';             -- endofpacket
			ff_tx_err     : in  std_logic                     := 'X';             -- error
			ff_tx_mod     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- empty
			ff_tx_rdy     : out std_logic;                                        -- ready
			ff_tx_sop     : in  std_logic                     := 'X';             -- startofpacket
			ff_tx_wren    : in  std_logic                     := 'X';             -- valid
			ff_tx_crc_fwd : in  std_logic                     := 'X';             -- ff_tx_crc_fwd
			ff_tx_septy   : out std_logic;                                        -- ff_tx_septy
			tx_ff_uflow   : out std_logic;                                        -- tx_ff_uflow
			ff_tx_a_full  : out std_logic;                                        -- ff_tx_a_full
			ff_tx_a_empty : out std_logic;                                        -- ff_tx_a_empty
			rx_err_stat   : out std_logic_vector(17 downto 0);                    -- rx_err_stat
			rx_frm_type   : out std_logic_vector(3 downto 0);                     -- rx_frm_type
			ff_rx_dsav    : out std_logic;                                        -- ff_rx_dsav
			ff_rx_a_full  : out std_logic;                                        -- ff_rx_a_full
			ff_rx_a_empty : out std_logic                                         -- ff_rx_a_empty
		);
	end component ethernet_setup_eth_tse_0;

	component ethernet_setup_jtaguart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component ethernet_setup_jtaguart_0;

	component ethernet_setup_nios2_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(16 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(16 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component ethernet_setup_nios2_0;

	component ethernet_setup_onchip_memory2_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component ethernet_setup_onchip_memory2_0;

	component ethernet_setup_sysid_qsys_0 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component ethernet_setup_sysid_qsys_0;

	component ethernet_setup_timer_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component ethernet_setup_timer_0;

	component ethernet_setup_mm_interconnect_0 is
		port (
			altpll_0_c1_clk                                            : in  std_logic                     := 'X';             -- clk
			clk_0_clk_clk                                              : in  std_logic                     := 'X';             -- clk
			altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			nios2_0_reset_reset_bridge_in_reset_reset                  : in  std_logic                     := 'X';             -- reset
			timer_0_reset_reset_bridge_in_reset_reset                  : in  std_logic                     := 'X';             -- reset
			nios2_0_data_master_address                                : in  std_logic_vector(16 downto 0) := (others => 'X'); -- address
			nios2_0_data_master_waitrequest                            : out std_logic;                                        -- waitrequest
			nios2_0_data_master_byteenable                             : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_0_data_master_read                                   : in  std_logic                     := 'X';             -- read
			nios2_0_data_master_readdata                               : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_0_data_master_readdatavalid                          : out std_logic;                                        -- readdatavalid
			nios2_0_data_master_write                                  : in  std_logic                     := 'X';             -- write
			nios2_0_data_master_writedata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_0_data_master_debugaccess                            : in  std_logic                     := 'X';             -- debugaccess
			nios2_0_instruction_master_address                         : in  std_logic_vector(16 downto 0) := (others => 'X'); -- address
			nios2_0_instruction_master_waitrequest                     : out std_logic;                                        -- waitrequest
			nios2_0_instruction_master_read                            : in  std_logic                     := 'X';             -- read
			nios2_0_instruction_master_readdata                        : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_0_instruction_master_readdatavalid                   : out std_logic;                                        -- readdatavalid
			altpll_0_pll_slave_address                                 : out std_logic_vector(1 downto 0);                     -- address
			altpll_0_pll_slave_write                                   : out std_logic;                                        -- write
			altpll_0_pll_slave_read                                    : out std_logic;                                        -- read
			altpll_0_pll_slave_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			altpll_0_pll_slave_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			eth_tse_0_control_port_address                             : out std_logic_vector(7 downto 0);                     -- address
			eth_tse_0_control_port_write                               : out std_logic;                                        -- write
			eth_tse_0_control_port_read                                : out std_logic;                                        -- read
			eth_tse_0_control_port_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			eth_tse_0_control_port_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			eth_tse_0_control_port_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			jtaguart_0_avalon_jtag_slave_address                       : out std_logic_vector(0 downto 0);                     -- address
			jtaguart_0_avalon_jtag_slave_write                         : out std_logic;                                        -- write
			jtaguart_0_avalon_jtag_slave_read                          : out std_logic;                                        -- read
			jtaguart_0_avalon_jtag_slave_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtaguart_0_avalon_jtag_slave_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			jtaguart_0_avalon_jtag_slave_waitrequest                   : in  std_logic                     := 'X';             -- waitrequest
			jtaguart_0_avalon_jtag_slave_chipselect                    : out std_logic;                                        -- chipselect
			nios2_0_debug_mem_slave_address                            : out std_logic_vector(8 downto 0);                     -- address
			nios2_0_debug_mem_slave_write                              : out std_logic;                                        -- write
			nios2_0_debug_mem_slave_read                               : out std_logic;                                        -- read
			nios2_0_debug_mem_slave_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_0_debug_mem_slave_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_0_debug_mem_slave_byteenable                         : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_0_debug_mem_slave_waitrequest                        : in  std_logic                     := 'X';             -- waitrequest
			nios2_0_debug_mem_slave_debugaccess                        : out std_logic;                                        -- debugaccess
			onchip_memory2_0_s1_address                                : out std_logic_vector(12 downto 0);                    -- address
			onchip_memory2_0_s1_write                                  : out std_logic;                                        -- write
			onchip_memory2_0_s1_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_0_s1_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_0_s1_byteenable                             : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_0_s1_chipselect                             : out std_logic;                                        -- chipselect
			onchip_memory2_0_s1_clken                                  : out std_logic;                                        -- clken
			sysid_qsys_0_control_slave_address                         : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_0_control_slave_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_address                                         : out std_logic_vector(2 downto 0);                     -- address
			timer_0_s1_write                                           : out std_logic;                                        -- write
			timer_0_s1_readdata                                        : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_writedata                                       : out std_logic_vector(15 downto 0);                    -- writedata
			timer_0_s1_chipselect                                      : out std_logic                                         -- chipselect
		);
	end component ethernet_setup_mm_interconnect_0;

	component ethernet_setup_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component ethernet_setup_irq_mapper;

	component ethernet_setup_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component ethernet_setup_rst_controller;

	component ethernet_setup_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component ethernet_setup_rst_controller_001;

	signal altpll_0_c0_clk                                                : std_logic;                     -- altpll_0:c0 -> [eth_tse_0:ff_rx_clk, eth_tse_0:ff_tx_clk, eth_tse_0:rx_clk, eth_tse_0:tx_clk]
	signal altpll_0_c1_clk                                                : std_logic;                     -- altpll_0:c1 -> [eth_tse_0:clk, irq_mapper:clk, jtaguart_0:clk, mm_interconnect_0:altpll_0_c1_clk, nios2_0:clk, onchip_memory2_0:clk, rst_controller_001:clk, rst_controller_002:clk, sysid_qsys_0:clock, timer_0:clk]
	signal nios2_0_data_master_readdata                                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_0_data_master_readdata -> nios2_0:d_readdata
	signal nios2_0_data_master_waitrequest                                : std_logic;                     -- mm_interconnect_0:nios2_0_data_master_waitrequest -> nios2_0:d_waitrequest
	signal nios2_0_data_master_debugaccess                                : std_logic;                     -- nios2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_0_data_master_debugaccess
	signal nios2_0_data_master_address                                    : std_logic_vector(16 downto 0); -- nios2_0:d_address -> mm_interconnect_0:nios2_0_data_master_address
	signal nios2_0_data_master_byteenable                                 : std_logic_vector(3 downto 0);  -- nios2_0:d_byteenable -> mm_interconnect_0:nios2_0_data_master_byteenable
	signal nios2_0_data_master_read                                       : std_logic;                     -- nios2_0:d_read -> mm_interconnect_0:nios2_0_data_master_read
	signal nios2_0_data_master_readdatavalid                              : std_logic;                     -- mm_interconnect_0:nios2_0_data_master_readdatavalid -> nios2_0:d_readdatavalid
	signal nios2_0_data_master_write                                      : std_logic;                     -- nios2_0:d_write -> mm_interconnect_0:nios2_0_data_master_write
	signal nios2_0_data_master_writedata                                  : std_logic_vector(31 downto 0); -- nios2_0:d_writedata -> mm_interconnect_0:nios2_0_data_master_writedata
	signal nios2_0_instruction_master_readdata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_0_instruction_master_readdata -> nios2_0:i_readdata
	signal nios2_0_instruction_master_waitrequest                         : std_logic;                     -- mm_interconnect_0:nios2_0_instruction_master_waitrequest -> nios2_0:i_waitrequest
	signal nios2_0_instruction_master_address                             : std_logic_vector(16 downto 0); -- nios2_0:i_address -> mm_interconnect_0:nios2_0_instruction_master_address
	signal nios2_0_instruction_master_read                                : std_logic;                     -- nios2_0:i_read -> mm_interconnect_0:nios2_0_instruction_master_read
	signal nios2_0_instruction_master_readdatavalid                       : std_logic;                     -- mm_interconnect_0:nios2_0_instruction_master_readdatavalid -> nios2_0:i_readdatavalid
	signal mm_interconnect_0_jtaguart_0_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtaguart_0_avalon_jtag_slave_chipselect -> jtaguart_0:av_chipselect
	signal mm_interconnect_0_jtaguart_0_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtaguart_0:av_readdata -> mm_interconnect_0:jtaguart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtaguart_0_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtaguart_0:av_waitrequest -> mm_interconnect_0:jtaguart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtaguart_0_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtaguart_0_avalon_jtag_slave_address -> jtaguart_0:av_address
	signal mm_interconnect_0_jtaguart_0_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtaguart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtaguart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtaguart_0_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtaguart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtaguart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtaguart_0_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtaguart_0_avalon_jtag_slave_writedata -> jtaguart_0:av_writedata
	signal mm_interconnect_0_eth_tse_0_control_port_readdata              : std_logic_vector(31 downto 0); -- eth_tse_0:reg_data_out -> mm_interconnect_0:eth_tse_0_control_port_readdata
	signal mm_interconnect_0_eth_tse_0_control_port_waitrequest           : std_logic;                     -- eth_tse_0:reg_busy -> mm_interconnect_0:eth_tse_0_control_port_waitrequest
	signal mm_interconnect_0_eth_tse_0_control_port_address               : std_logic_vector(7 downto 0);  -- mm_interconnect_0:eth_tse_0_control_port_address -> eth_tse_0:reg_addr
	signal mm_interconnect_0_eth_tse_0_control_port_read                  : std_logic;                     -- mm_interconnect_0:eth_tse_0_control_port_read -> eth_tse_0:reg_rd
	signal mm_interconnect_0_eth_tse_0_control_port_write                 : std_logic;                     -- mm_interconnect_0:eth_tse_0_control_port_write -> eth_tse_0:reg_wr
	signal mm_interconnect_0_eth_tse_0_control_port_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:eth_tse_0_control_port_writedata -> eth_tse_0:reg_data_in
	signal mm_interconnect_0_sysid_qsys_0_control_slave_readdata          : std_logic_vector(31 downto 0); -- sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_address           : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	signal mm_interconnect_0_nios2_0_debug_mem_slave_readdata             : std_logic_vector(31 downto 0); -- nios2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_0_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_0_debug_mem_slave_waitrequest          : std_logic;                     -- nios2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_0_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_0_debug_mem_slave_debugaccess          : std_logic;                     -- mm_interconnect_0:nios2_0_debug_mem_slave_debugaccess -> nios2_0:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_0_debug_mem_slave_address              : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_0_debug_mem_slave_address -> nios2_0:debug_mem_slave_address
	signal mm_interconnect_0_nios2_0_debug_mem_slave_read                 : std_logic;                     -- mm_interconnect_0:nios2_0_debug_mem_slave_read -> nios2_0:debug_mem_slave_read
	signal mm_interconnect_0_nios2_0_debug_mem_slave_byteenable           : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_0_debug_mem_slave_byteenable -> nios2_0:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_0_debug_mem_slave_write                : std_logic;                     -- mm_interconnect_0:nios2_0_debug_mem_slave_write -> nios2_0:debug_mem_slave_write
	signal mm_interconnect_0_nios2_0_debug_mem_slave_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_0_debug_mem_slave_writedata -> nios2_0:debug_mem_slave_writedata
	signal mm_interconnect_0_altpll_0_pll_slave_readdata                  : std_logic_vector(31 downto 0); -- altpll_0:readdata -> mm_interconnect_0:altpll_0_pll_slave_readdata
	signal mm_interconnect_0_altpll_0_pll_slave_address                   : std_logic_vector(1 downto 0);  -- mm_interconnect_0:altpll_0_pll_slave_address -> altpll_0:address
	signal mm_interconnect_0_altpll_0_pll_slave_read                      : std_logic;                     -- mm_interconnect_0:altpll_0_pll_slave_read -> altpll_0:read
	signal mm_interconnect_0_altpll_0_pll_slave_write                     : std_logic;                     -- mm_interconnect_0:altpll_0_pll_slave_write -> altpll_0:write
	signal mm_interconnect_0_altpll_0_pll_slave_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:altpll_0_pll_slave_writedata -> altpll_0:writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_chipselect               : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	signal mm_interconnect_0_onchip_memory2_0_s1_readdata                 : std_logic_vector(31 downto 0); -- onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	signal mm_interconnect_0_onchip_memory2_0_s1_address                  : std_logic_vector(12 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	signal mm_interconnect_0_onchip_memory2_0_s1_byteenable               : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	signal mm_interconnect_0_onchip_memory2_0_s1_write                    : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	signal mm_interconnect_0_onchip_memory2_0_s1_writedata                : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_clken                    : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	signal mm_interconnect_0_timer_0_s1_chipselect                        : std_logic;                     -- mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	signal mm_interconnect_0_timer_0_s1_readdata                          : std_logic_vector(15 downto 0); -- timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	signal mm_interconnect_0_timer_0_s1_address                           : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_0_s1_address -> timer_0:address
	signal mm_interconnect_0_timer_0_s1_write                             : std_logic;                     -- mm_interconnect_0:timer_0_s1_write -> mm_interconnect_0_timer_0_s1_write:in
	signal mm_interconnect_0_timer_0_s1_writedata                         : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	signal irq_mapper_receiver0_irq                                       : std_logic;                     -- jtaguart_0:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                       : std_logic;                     -- timer_0:irq -> irq_mapper:receiver1_irq
	signal nios2_0_irq_irq                                                : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_0:irq
	signal rst_controller_reset_out_reset                                 : std_logic;                     -- rst_controller:reset_out -> [altpll_0:reset, mm_interconnect_0:altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset]
	signal rst_controller_001_reset_out_reset                             : std_logic;                     -- rst_controller_001:reset_out -> [eth_tse_0:reset, irq_mapper:reset, mm_interconnect_0:nios2_0_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_controller_001_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_001_reset_out_reset_req                         : std_logic;                     -- rst_controller_001:reset_req -> [nios2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	signal nios2_0_debug_reset_request_reset                              : std_logic;                     -- nios2_0:debug_reset_request -> rst_controller_001:reset_in1
	signal rst_controller_002_reset_out_reset                             : std_logic;                     -- rst_controller_002:reset_out -> [mm_interconnect_0:timer_0_reset_reset_bridge_in_reset_reset, rst_controller_002_reset_out_reset:in]
	signal reset_reset_n_ports_inv                                        : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0]
	signal mm_interconnect_0_jtaguart_0_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtaguart_0_avalon_jtag_slave_read:inv -> jtaguart_0:av_read_n
	signal mm_interconnect_0_jtaguart_0_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtaguart_0_avalon_jtag_slave_write:inv -> jtaguart_0:av_write_n
	signal mm_interconnect_0_timer_0_s1_write_ports_inv                   : std_logic;                     -- mm_interconnect_0_timer_0_s1_write:inv -> timer_0:write_n
	signal rst_controller_001_reset_out_reset_ports_inv                   : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [jtaguart_0:rst_n, nios2_0:reset_n, sysid_qsys_0:reset_n]
	signal rst_controller_002_reset_out_reset_ports_inv                   : std_logic;                     -- rst_controller_002_reset_out_reset:inv -> timer_0:reset_n

begin

	altpll_0 : component ethernet_setup_altpll_0
		port map (
			clk                => clk_clk,                                        --       inclk_interface.clk
			reset              => rst_controller_reset_out_reset,                 -- inclk_interface_reset.reset
			read               => mm_interconnect_0_altpll_0_pll_slave_read,      --             pll_slave.read
			write              => mm_interconnect_0_altpll_0_pll_slave_write,     --                      .write
			address            => mm_interconnect_0_altpll_0_pll_slave_address,   --                      .address
			readdata           => mm_interconnect_0_altpll_0_pll_slave_readdata,  --                      .readdata
			writedata          => mm_interconnect_0_altpll_0_pll_slave_writedata, --                      .writedata
			c0                 => altpll_0_c0_clk,                                --                    c0.clk
			c1                 => altpll_0_c1_clk,                                --                    c1.clk
			c2                 => altpll_0_c2_clk,                                --                    c2.clk
			areset             => altpll_0_areset_conduit_export,                 --        areset_conduit.export
			locked             => altpll_0_locked_conduit_export,                 --        locked_conduit.export
			scandone           => open,                                           --           (terminated)
			scandataout        => open,                                           --           (terminated)
			c3                 => open,                                           --           (terminated)
			c4                 => open,                                           --           (terminated)
			phasedone          => open,                                           --           (terminated)
			phasecounterselect => "000",                                          --           (terminated)
			phaseupdown        => '0',                                            --           (terminated)
			phasestep          => '0',                                            --           (terminated)
			scanclk            => '0',                                            --           (terminated)
			scanclkena         => '0',                                            --           (terminated)
			scandata           => '0',                                            --           (terminated)
			configupdate       => '0'                                             --           (terminated)
		);

	eth_tse_0 : component ethernet_setup_eth_tse_0
		port map (
			clk           => altpll_0_c1_clk,                                      -- control_port_clock_connection.clk
			reset         => rst_controller_001_reset_out_reset,                   --              reset_connection.reset
			reg_addr      => mm_interconnect_0_eth_tse_0_control_port_address,     --                  control_port.address
			reg_data_out  => mm_interconnect_0_eth_tse_0_control_port_readdata,    --                              .readdata
			reg_rd        => mm_interconnect_0_eth_tse_0_control_port_read,        --                              .read
			reg_data_in   => mm_interconnect_0_eth_tse_0_control_port_writedata,   --                              .writedata
			reg_wr        => mm_interconnect_0_eth_tse_0_control_port_write,       --                              .write
			reg_busy      => mm_interconnect_0_eth_tse_0_control_port_waitrequest, --                              .waitrequest
			tx_clk        => altpll_0_c0_clk,                                      --   pcs_mac_tx_clock_connection.clk
			rx_clk        => altpll_0_c0_clk,                                      --   pcs_mac_rx_clock_connection.clk
			set_10        => eth_tse_0_mac_status_connection_set_10,               --         mac_status_connection.set_10
			set_1000      => eth_tse_0_mac_status_connection_set_1000,             --                              .set_1000
			eth_mode      => eth_tse_0_mac_status_connection_eth_mode,             --                              .eth_mode
			ena_10        => eth_tse_0_mac_status_connection_ena_10,               --                              .ena_10
			rgmii_in      => eth_tse_0_mac_rgmii_connection_rgmii_in,              --          mac_rgmii_connection.rgmii_in
			rgmii_out     => eth_tse_0_mac_rgmii_connection_rgmii_out,             --                              .rgmii_out
			rx_control    => eth_tse_0_mac_rgmii_connection_rx_control,            --                              .rx_control
			tx_control    => eth_tse_0_mac_rgmii_connection_tx_control,            --                              .tx_control
			ff_rx_clk     => altpll_0_c0_clk,                                      --      receive_clock_connection.clk
			ff_tx_clk     => altpll_0_c0_clk,                                      --     transmit_clock_connection.clk
			ff_rx_data    => eth_tse_0_receive_data,                               --                       receive.data
			ff_rx_eop     => eth_tse_0_receive_endofpacket,                        --                              .endofpacket
			rx_err        => eth_tse_0_receive_error,                              --                              .error
			ff_rx_mod     => eth_tse_0_receive_empty,                              --                              .empty
			ff_rx_rdy     => eth_tse_0_receive_ready,                              --                              .ready
			ff_rx_sop     => eth_tse_0_receive_startofpacket,                      --                              .startofpacket
			ff_rx_dval    => eth_tse_0_receive_valid,                              --                              .valid
			ff_tx_data    => eth_tse_0_transmit_data,                              --                      transmit.data
			ff_tx_eop     => eth_tse_0_transmit_endofpacket,                       --                              .endofpacket
			ff_tx_err     => eth_tse_0_transmit_error,                             --                              .error
			ff_tx_mod     => eth_tse_0_transmit_empty,                             --                              .empty
			ff_tx_rdy     => eth_tse_0_transmit_ready,                             --                              .ready
			ff_tx_sop     => eth_tse_0_transmit_startofpacket,                     --                              .startofpacket
			ff_tx_wren    => eth_tse_0_transmit_valid,                             --                              .valid
			ff_tx_crc_fwd => eth_tse_0_mac_misc_connection_ff_tx_crc_fwd,          --           mac_misc_connection.ff_tx_crc_fwd
			ff_tx_septy   => eth_tse_0_mac_misc_connection_ff_tx_septy,            --                              .ff_tx_septy
			tx_ff_uflow   => eth_tse_0_mac_misc_connection_tx_ff_uflow,            --                              .tx_ff_uflow
			ff_tx_a_full  => eth_tse_0_mac_misc_connection_ff_tx_a_full,           --                              .ff_tx_a_full
			ff_tx_a_empty => eth_tse_0_mac_misc_connection_ff_tx_a_empty,          --                              .ff_tx_a_empty
			rx_err_stat   => eth_tse_0_mac_misc_connection_rx_err_stat,            --                              .rx_err_stat
			rx_frm_type   => eth_tse_0_mac_misc_connection_rx_frm_type,            --                              .rx_frm_type
			ff_rx_dsav    => eth_tse_0_mac_misc_connection_ff_rx_dsav,             --                              .ff_rx_dsav
			ff_rx_a_full  => eth_tse_0_mac_misc_connection_ff_rx_a_full,           --                              .ff_rx_a_full
			ff_rx_a_empty => eth_tse_0_mac_misc_connection_ff_rx_a_empty           --                              .ff_rx_a_empty
		);

	jtaguart_0 : component ethernet_setup_jtaguart_0
		port map (
			clk            => altpll_0_c1_clk,                                                --               clk.clk
			rst_n          => rst_controller_001_reset_out_reset_ports_inv,                   --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtaguart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtaguart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtaguart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtaguart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtaguart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtaguart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtaguart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                        --               irq.irq
		);

	nios2_0 : component ethernet_setup_nios2_0
		port map (
			clk                                 => altpll_0_c1_clk,                                       --                       clk.clk
			reset_n                             => rst_controller_001_reset_out_reset_ports_inv,          --                     reset.reset_n
			reset_req                           => rst_controller_001_reset_out_reset_req,                --                          .reset_req
			d_address                           => nios2_0_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_0_data_master_read,                              --                          .read
			d_readdata                          => nios2_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_0_data_master_write,                             --                          .write
			d_writedata                         => nios2_0_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => nios2_0_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => nios2_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_0_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_0_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => nios2_0_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => nios2_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_0_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                   -- custom_instruction_master.readra
		);

	onchip_memory2_0 : component ethernet_setup_onchip_memory2_0
		port map (
			clk        => altpll_0_c1_clk,                                  --   clk1.clk
			address    => mm_interconnect_0_onchip_memory2_0_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory2_0_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory2_0_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory2_0_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory2_0_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory2_0_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory2_0_s1_byteenable, --       .byteenable
			reset      => rst_controller_001_reset_out_reset,               -- reset1.reset
			reset_req  => rst_controller_001_reset_out_reset_req,           --       .reset_req
			freeze     => '0'                                               -- (terminated)
		);

	sysid_qsys_0 : component ethernet_setup_sysid_qsys_0
		port map (
			clock    => altpll_0_c1_clk,                                         --           clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv,            --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_0_control_slave_address(0)  --              .address
		);

	timer_0 : component ethernet_setup_timer_0
		port map (
			clk        => altpll_0_c1_clk,                              --   clk.clk
			reset_n    => rst_controller_002_reset_out_reset_ports_inv, -- reset.reset_n
			address    => mm_interconnect_0_timer_0_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_0_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_0_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_0_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_0_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver1_irq                      --   irq.irq
		);

	mm_interconnect_0 : component ethernet_setup_mm_interconnect_0
		port map (
			altpll_0_c1_clk                                            => altpll_0_c1_clk,                                            --                                          altpll_0_c1.clk
			clk_0_clk_clk                                              => clk_clk,                                                    --                                            clk_0_clk.clk
			altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                             -- altpll_0_inclk_interface_reset_reset_bridge_in_reset.reset
			nios2_0_reset_reset_bridge_in_reset_reset                  => rst_controller_001_reset_out_reset,                         --                  nios2_0_reset_reset_bridge_in_reset.reset
			timer_0_reset_reset_bridge_in_reset_reset                  => rst_controller_002_reset_out_reset,                         --                  timer_0_reset_reset_bridge_in_reset.reset
			nios2_0_data_master_address                                => nios2_0_data_master_address,                                --                                  nios2_0_data_master.address
			nios2_0_data_master_waitrequest                            => nios2_0_data_master_waitrequest,                            --                                                     .waitrequest
			nios2_0_data_master_byteenable                             => nios2_0_data_master_byteenable,                             --                                                     .byteenable
			nios2_0_data_master_read                                   => nios2_0_data_master_read,                                   --                                                     .read
			nios2_0_data_master_readdata                               => nios2_0_data_master_readdata,                               --                                                     .readdata
			nios2_0_data_master_readdatavalid                          => nios2_0_data_master_readdatavalid,                          --                                                     .readdatavalid
			nios2_0_data_master_write                                  => nios2_0_data_master_write,                                  --                                                     .write
			nios2_0_data_master_writedata                              => nios2_0_data_master_writedata,                              --                                                     .writedata
			nios2_0_data_master_debugaccess                            => nios2_0_data_master_debugaccess,                            --                                                     .debugaccess
			nios2_0_instruction_master_address                         => nios2_0_instruction_master_address,                         --                           nios2_0_instruction_master.address
			nios2_0_instruction_master_waitrequest                     => nios2_0_instruction_master_waitrequest,                     --                                                     .waitrequest
			nios2_0_instruction_master_read                            => nios2_0_instruction_master_read,                            --                                                     .read
			nios2_0_instruction_master_readdata                        => nios2_0_instruction_master_readdata,                        --                                                     .readdata
			nios2_0_instruction_master_readdatavalid                   => nios2_0_instruction_master_readdatavalid,                   --                                                     .readdatavalid
			altpll_0_pll_slave_address                                 => mm_interconnect_0_altpll_0_pll_slave_address,               --                                   altpll_0_pll_slave.address
			altpll_0_pll_slave_write                                   => mm_interconnect_0_altpll_0_pll_slave_write,                 --                                                     .write
			altpll_0_pll_slave_read                                    => mm_interconnect_0_altpll_0_pll_slave_read,                  --                                                     .read
			altpll_0_pll_slave_readdata                                => mm_interconnect_0_altpll_0_pll_slave_readdata,              --                                                     .readdata
			altpll_0_pll_slave_writedata                               => mm_interconnect_0_altpll_0_pll_slave_writedata,             --                                                     .writedata
			eth_tse_0_control_port_address                             => mm_interconnect_0_eth_tse_0_control_port_address,           --                               eth_tse_0_control_port.address
			eth_tse_0_control_port_write                               => mm_interconnect_0_eth_tse_0_control_port_write,             --                                                     .write
			eth_tse_0_control_port_read                                => mm_interconnect_0_eth_tse_0_control_port_read,              --                                                     .read
			eth_tse_0_control_port_readdata                            => mm_interconnect_0_eth_tse_0_control_port_readdata,          --                                                     .readdata
			eth_tse_0_control_port_writedata                           => mm_interconnect_0_eth_tse_0_control_port_writedata,         --                                                     .writedata
			eth_tse_0_control_port_waitrequest                         => mm_interconnect_0_eth_tse_0_control_port_waitrequest,       --                                                     .waitrequest
			jtaguart_0_avalon_jtag_slave_address                       => mm_interconnect_0_jtaguart_0_avalon_jtag_slave_address,     --                         jtaguart_0_avalon_jtag_slave.address
			jtaguart_0_avalon_jtag_slave_write                         => mm_interconnect_0_jtaguart_0_avalon_jtag_slave_write,       --                                                     .write
			jtaguart_0_avalon_jtag_slave_read                          => mm_interconnect_0_jtaguart_0_avalon_jtag_slave_read,        --                                                     .read
			jtaguart_0_avalon_jtag_slave_readdata                      => mm_interconnect_0_jtaguart_0_avalon_jtag_slave_readdata,    --                                                     .readdata
			jtaguart_0_avalon_jtag_slave_writedata                     => mm_interconnect_0_jtaguart_0_avalon_jtag_slave_writedata,   --                                                     .writedata
			jtaguart_0_avalon_jtag_slave_waitrequest                   => mm_interconnect_0_jtaguart_0_avalon_jtag_slave_waitrequest, --                                                     .waitrequest
			jtaguart_0_avalon_jtag_slave_chipselect                    => mm_interconnect_0_jtaguart_0_avalon_jtag_slave_chipselect,  --                                                     .chipselect
			nios2_0_debug_mem_slave_address                            => mm_interconnect_0_nios2_0_debug_mem_slave_address,          --                              nios2_0_debug_mem_slave.address
			nios2_0_debug_mem_slave_write                              => mm_interconnect_0_nios2_0_debug_mem_slave_write,            --                                                     .write
			nios2_0_debug_mem_slave_read                               => mm_interconnect_0_nios2_0_debug_mem_slave_read,             --                                                     .read
			nios2_0_debug_mem_slave_readdata                           => mm_interconnect_0_nios2_0_debug_mem_slave_readdata,         --                                                     .readdata
			nios2_0_debug_mem_slave_writedata                          => mm_interconnect_0_nios2_0_debug_mem_slave_writedata,        --                                                     .writedata
			nios2_0_debug_mem_slave_byteenable                         => mm_interconnect_0_nios2_0_debug_mem_slave_byteenable,       --                                                     .byteenable
			nios2_0_debug_mem_slave_waitrequest                        => mm_interconnect_0_nios2_0_debug_mem_slave_waitrequest,      --                                                     .waitrequest
			nios2_0_debug_mem_slave_debugaccess                        => mm_interconnect_0_nios2_0_debug_mem_slave_debugaccess,      --                                                     .debugaccess
			onchip_memory2_0_s1_address                                => mm_interconnect_0_onchip_memory2_0_s1_address,              --                                  onchip_memory2_0_s1.address
			onchip_memory2_0_s1_write                                  => mm_interconnect_0_onchip_memory2_0_s1_write,                --                                                     .write
			onchip_memory2_0_s1_readdata                               => mm_interconnect_0_onchip_memory2_0_s1_readdata,             --                                                     .readdata
			onchip_memory2_0_s1_writedata                              => mm_interconnect_0_onchip_memory2_0_s1_writedata,            --                                                     .writedata
			onchip_memory2_0_s1_byteenable                             => mm_interconnect_0_onchip_memory2_0_s1_byteenable,           --                                                     .byteenable
			onchip_memory2_0_s1_chipselect                             => mm_interconnect_0_onchip_memory2_0_s1_chipselect,           --                                                     .chipselect
			onchip_memory2_0_s1_clken                                  => mm_interconnect_0_onchip_memory2_0_s1_clken,                --                                                     .clken
			sysid_qsys_0_control_slave_address                         => mm_interconnect_0_sysid_qsys_0_control_slave_address,       --                           sysid_qsys_0_control_slave.address
			sysid_qsys_0_control_slave_readdata                        => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,      --                                                     .readdata
			timer_0_s1_address                                         => mm_interconnect_0_timer_0_s1_address,                       --                                           timer_0_s1.address
			timer_0_s1_write                                           => mm_interconnect_0_timer_0_s1_write,                         --                                                     .write
			timer_0_s1_readdata                                        => mm_interconnect_0_timer_0_s1_readdata,                      --                                                     .readdata
			timer_0_s1_writedata                                       => mm_interconnect_0_timer_0_s1_writedata,                     --                                                     .writedata
			timer_0_s1_chipselect                                      => mm_interconnect_0_timer_0_s1_chipselect                     --                                                     .chipselect
		);

	irq_mapper : component ethernet_setup_irq_mapper
		port map (
			clk           => altpll_0_c1_clk,                    --       clk.clk
			reset         => rst_controller_001_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			sender_irq    => nios2_0_irq_irq                     --    sender.irq
		);

	rst_controller : component ethernet_setup_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component ethernet_setup_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			reset_in1      => nios2_0_debug_reset_request_reset,      -- reset_in1.reset
			clk            => altpll_0_c1_clk,                        --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_001_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_002 : component ethernet_setup_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => altpll_0_c1_clk,                    --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtaguart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtaguart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtaguart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtaguart_0_avalon_jtag_slave_write;

	mm_interconnect_0_timer_0_s1_write_ports_inv <= not mm_interconnect_0_timer_0_s1_write;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

end architecture rtl; -- of ethernet_setup
