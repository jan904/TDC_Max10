-- Channel for signal detection. This module detects the signal and encodes its timing information.

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_arith.ALL;

ENTITY channel IS
    GENERIC (
        carry4_count : INTEGER := 72;                                       -- carry4_count * 4: Number of bins in the delay line
        n_output_bits : INTEGER := 9                                        -- Number of bits for fine timestamp
    );
    PORT (  
        clk : IN STD_LOGIC;                                                 -- Clock Input               
        signal_in : IN STD_LOGIC;                                           -- Input signal which is to be detected
        start_reset : IN STD_LOGIC;                                         -- Reset signal after start of the FPGA. Generated by handle_start
        channel_written : IN STD_LOGIC;                                     -- Signal to indicate that the output of this channel has been written to the FIFO
        signal_out : OUT STD_LOGIC_VECTOR(n_output_bits - 1 DOWNTO 0);      -- Fine timestamp output
        wr_en_out : OUT STD_LOGIC                                           -- Write enable: Indicates that the output of this channel is ready to be written to the FIFO
    );
END ENTITY channel;


ARCHITECTURE rtl OF channel IS

    SIGNAL reset_after_signal : STD_LOGIC;
    SIGNAL busy : STD_LOGIC;
    SIGNAL wr_en : STD_LOGIC;
    SIGNAL therm_code : STD_LOGIC_VECTOR(carry4_count * 4 - 1 DOWNTO 0);
    SIGNAL bin_output : STD_LOGIC_VECTOR(n_output_bits - 1 DOWNTO 0);

    COMPONENT delay_line IS
        GENERIC (
            stages : POSITIVE
        );
        PORT (
            reset : IN STD_LOGIC;
            trigger : IN STD_LOGIC;
            clock : IN STD_LOGIC;
            signal_running : IN STD_LOGIC;
            therm_code : OUT STD_LOGIC_VECTOR(stages - 1 DOWNTO 0)
        );
    END COMPONENT delay_line;

    COMPONENT encoder IS
        GENERIC (
            n_bits_bin : POSITIVE;
            n_bits_therm : POSITIVE
        );
        PORT (
            clk : IN STD_LOGIC;
            thermometer : IN STD_LOGIC_VECTOR((n_bits_therm - 1) DOWNTO 0);
            count_bin : OUT STD_LOGIC_VECTOR(n_bits_bin - 1 DOWNTO 0)
        );
    END COMPONENT encoder;

    COMPONENT detect_signal IS
        GENERIC (
            stages : POSITIVE;
            n_output_bits : POSITIVE
        );
        PORT (
            clock : IN STD_LOGIC;
            start : IN STD_LOGIC;
            signal_in : IN STD_LOGIC;
            written : IN STD_LOGIC;
            signal_running : OUT STD_LOGIC;
            reset : OUT STD_LOGIC;
            wrt : OUT STD_LOGIC
        );
    END COMPONENT detect_signal;

BEGIN

    -- Actual delay line of delay elements
    delay_line_inst : delay_line
    GENERIC MAP(
        stages => carry4_count * 4
    )
    PORT MAP(
        reset => reset_after_signal,
        signal_running => busy,
        trigger => signal_in,
        clock => clk,
        therm_code => therm_code
    );
	 
    -- Detect incoming signal and handle status signals
    detect_signal_inst : detect_signal
    GENERIC MAP(
        stages => carry4_count * 4,
        n_output_bits => n_output_bits
    )
    PORT MAP(
        clock => clk,
        start => start_reset,
        signal_in => signal_in,
        written => channel_written,
        signal_running => busy,
        reset => reset_after_signal,
        wrt => wr_en_out
    );
	 
    -- Encode the thermometer code to binary
    encoder_inst : encoder
    GENERIC MAP(
        n_bits_bin => n_output_bits,
        n_bits_therm => 4 * carry4_count
    )
    PORT MAP(
        clk => clk,
        thermometer => therm_code,
        count_bin => bin_output
    );

    -- Output the fine timestamp
    signal_out <= bin_output;
        
END ARCHITECTURE rtl;